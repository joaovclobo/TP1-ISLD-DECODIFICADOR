module testeTp_tb;
reg [0:4] inp_teste;
wire [0:6] out_saida;

tp1isl uut (.entrada(inp_teste), .saida(out_saida));

initial begin
        $dumpfile("testeTp_tb.vcd");
        $dumpvars(0, testeTp_tb);
        $display("Comeco");

        #0 inp_teste = 5'b00000;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00001;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00010;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00011;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00100;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00101;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00110;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b00111;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01000;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01001;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01010;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01011;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01100;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01101;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01110;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b01111;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10000;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10001;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10010;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10011;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10100;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10101;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10110;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b10111;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11000;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11001;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11010;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11011;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11100;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11101;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11110;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #1 inp_teste = 5'b11111;
        $monitor("Entrada %b - Saida = %b", inp_teste, out_saida);
        #10 $stop;
        $display("Fim");
    end

endmodule